module tb ();
    reg clk;
    reg rstn;
    reg [15:0] bus;

  	datapath datapath1 (clk, rstn, bus);

    always #10 clk = ~clk;

    initial begin
      $dumpfile("dump.vcd");
      $dumpvars(0, tb);
    end


    initial begin
        clk = 0;
        rstn = 0;
      
        #20 rstn = 1;
    end

endmodule